real x [] = {
  1.10168563e+00,  1.38191166e+00,  1.29029608e+00,  1.05666263e+00,
  9.44225451e-01,  9.57986882e-01,  1.04630625e+00,  1.24103669e+00,
  1.44362822e+00,  1.38745155e+00,  1.03788056e+00,  7.75615544e-01,
  9.17805051e-01,  1.25377026e+00,  1.34262046e+00,  1.11761007e+00,
  8.80060491e-01,  8.01251778e-01,  7.82138913e-01,  7.71163204e-01,
  8.50151069e-01,  9.51564312e-01,  8.43666135e-01,  5.26837790e-01,
  3.34413249e-01,  4.60870481e-01,  6.60838912e-01,  6.31580228e-01,
  4.50306429e-01,  3.69054654e-01,  3.83036554e-01,  3.22866993e-01,
  2.34771114e-01,  3.09903368e-01,  4.88555652e-01,  4.94872306e-01,
  2.90170885e-01,  1.54792529e-01,  2.41699208e-01,  3.67060794e-01,
  3.67011578e-01,  3.52018911e-01,  4.22715296e-01,  4.22505237e-01,
  2.30924392e-01,  6.92671027e-02,  1.99402134e-01,  4.72317213e-01,
  5.11177191e-01,  2.62295942e-01,  3.17920701e-02,  4.35686085e-03,
  6.07462451e-02,  9.20818618e-02,  1.47698803e-01,  1.82786096e-01,
  4.17554112e-03, -3.60161193e-01, -5.43036481e-01, -3.30322882e-01,
 -3.10702896e-02, -7.89812886e-02, -4.44599871e-01, -7.39927603e-01,
 -7.72670233e-01, -6.76100854e-01, -5.76326523e-01, -4.84232970e-01,
 -5.01278126e-01, -7.62600670e-01, -1.10297157e+00, -1.12822054e+00,
 -7.68516036e-01, -4.58581970e-01, -5.70402768e-01, -9.25409361e-01,
 -1.10167650e+00, -9.98151934e-01, -8.18471327e-01, -6.82846507e-01,
 -5.84171074e-01, -6.09024981e-01, -8.39189875e-01, -1.06629994e+00,
 -9.65260886e-01, -5.96181604e-01, -3.99039690e-01, -5.91749772e-01,
 -8.86291631e-01, -9.45660659e-01, -8.22643699e-01, -7.41904480e-01,
 -7.20442206e-01, -6.77700826e-01, -7.07673975e-01, -9.16455200e-01,
 -1.12344019e+00, -1.06484800e+00, -8.32559680e-01, -7.75322055e-01,
 -9.74166119e-01, -1.15180838e+00, -1.14253457e+00, -1.10739966e+00,
 -1.17324544e+00, -1.19454037e+00, -1.06685594e+00, -9.85445284e-01,
 -1.13310647e+00, -1.33366307e+00, -1.30651078e+00, -1.10492217e+00,
 -9.97136728e-01, -1.02827509e+00, -1.02649315e+00, -9.75567758e-01,
 -1.02452668e+00, -1.12269355e+00, -1.01414213e+00, -6.89533517e-01,
 -5.01125046e-01, -6.58212204e-01, -8.98661577e-01, -8.76706068e-01,
 -6.33424086e-01, -4.37234862e-01, -3.68218495e-01, -3.46363592e-01,
 -4.01541400e-01, -5.79299038e-01, -6.79987056e-01, -4.59654445e-01,
 -7.84719499e-02,  1.22623524e-02, -3.04275466e-01, -6.27772770e-01,
 -5.98755735e-01, -3.34475208e-01, -1.49043724e-01, -1.27889994e-01,
 -1.98291745e-01, -3.63510191e-01, -5.81452831e-01, -6.09145302e-01,
 -3.02603705e-01,  4.43860658e-02,  7.25887135e-03, -3.67025504e-01,
 -6.01439901e-01, -4.40419019e-01, -1.25917883e-01,  3.50624550e-02,
  3.92751141e-02, -3.07175137e-03, -9.95560313e-02, -2.07904652e-01,
 -1.16300255e-01,  2.36885149e-01,  5.31641901e-01,  4.54743453e-01,
  1.74539639e-01,  1.16339456e-01,  3.62986024e-01,  6.10749546e-01,
  6.73872678e-01,  6.75097783e-01,  7.07827800e-01,  6.73207027e-01,
  5.68614863e-01,  6.05157873e-01,  8.50254713e-01,  1.03190328e+00,
  9.27826301e-01,  7.18797067e-01,  6.97472567e-01,  8.22020358e-01,
  8.56167381e-01,  8.00243003e-01,  8.38523930e-01,  9.37979388e-01,
  8.70544915e-01,  6.45208028e-01,  5.58961785e-01,  7.30252461e-01,
  9.05261245e-01,  8.65084489e-01,  7.31351304e-01,  6.89611265e-01,
  6.85037865e-01,  6.26191445e-01,  6.46149718e-01,  8.62053804e-01,
  1.05553885e+00,  9.37152439e-01,  6.33893653e-01,  5.61181787e-01,
  8.29465099e-01,  1.11639238e+00,  1.16132230e+00,  1.05707028e+00,
  9.69901751e-01,  9.00345235e-01,  8.69445225e-01,  1.02701240e+00,
  1.34826500e+00,  1.48761373e+00,  1.22187035e+00,  8.48298497e-01,
  8.28177007e-01,  1.15856707e+00,  1.41913905e+00,  1.36781530e+00,
  1.15537996e+00,  9.73822096e-01,  8.47271381e-01,  8.19558000e-01,
  9.90696203e-01,  1.23251918e+00,  1.19274289e+00,  7.87461668e-01,
  4.22354001e-01,  4.78397151e-01,  7.93268235e-01,  9.25593481e-01,
  7.57120612e-01,  5.25176411e-01,  3.88208474e-01,  3.08433495e-01,
  3.08051243e-01,  4.70872666e-01,  6.57791619e-01,  5.76054786e-01,
  2.38401223e-01,  3.59039151e-02,  1.98922078e-01,  4.70906647e-01,
  5.13415730e-01,  3.72131341e-01,  2.90997854e-01,  2.90876504e-01,
  2.44204087e-01,  2.08549418e-01,  3.34207349e-01,  5.13645740e-01,
  4.77516671e-01,  2.39954385e-01,  1.11346495e-01,  2.16843017e-01,
  3.28594879e-01,  2.76169850e-01,  1.99511077e-01,  2.27320329e-01,
  2.08488652e-01,  7.57506014e-03, -1.81275954e-01, -1.15757034e-01,
  7.23091231e-02,  5.69469770e-02, -1.86081274e-01, -3.87382350e-01,
 -4.28844913e-01, -4.44496946e-01, -4.85415695e-01, -4.39312105e-01,
 -3.50600374e-01, -4.66259129e-01, -8.08593977e-01, -1.01748101e+00,
 -8.41967989e-01, -5.35877878e-01, -5.03635650e-01, -7.50906323e-01,
 -9.69734007e-01, -1.01104022e+00, -9.58513773e-01, -8.45230138e-01,
 -6.50115561e-01, -5.37630582e-01, -7.28803003e-01, -1.08189942e+00,
 -1.15385587e+00, -8.06456440e-01, -4.41423215e-01, -4.57675530e-01,
 -7.48061563e-01, -9.47915188e-01, -9.36365636e-01, -8.28159517e-01,
 -6.76938938e-01, -5.07015305e-01, -4.99041318e-01, -7.86563296e-01,
 -1.12194859e+00, -1.10208216e+00, -7.47219060e-01, -5.18825063e-01,
 -6.89284681e-01, -1.01552593e+00, -1.15966504e+00, -1.11971197e+00,
 -1.05676254e+00, -9.84248350e-01, -8.88243028e-01, -9.25123529e-01,
 -1.18731242e+00, -1.42586092e+00, -1.33599473e+00, -1.03301621e+00,
 -9.14072842e-01, -1.08321874e+00, -1.25221744e+00, -1.22814971e+00,
 -1.14703012e+00, -1.13328401e+00, -1.07315455e+00, -9.01551158e-01,
 -8.11873578e-01, -9.39967936e-01, -1.07698753e+00, -9.69740591e-01,
 -7.24633724e-01, -6.20867804e-01, -6.63469090e-01, -6.43808971e-01,
 -5.51590021e-01, -5.68605361e-01, -6.69431351e-01, -6.00146496e-01,
 -3.28610366e-01, -1.69429968e-01, -3.12845699e-01, -5.28727778e-01,
 -5.31227338e-01, -3.77645630e-01, -2.78422939e-01, -2.43535833e-01,
 -1.92237154e-01, -2.21051059e-01, -4.32272976e-01, -6.17842567e-01,
 -4.77896483e-01, -1.21340140e-01,  1.00337395e-02, -2.41571968e-01,
 -5.41500644e-01, -5.61111188e-01, -3.69927171e-01, -1.93387002e-01,
 -8.40998383e-02, -3.52644901e-02, -1.44004916e-01, -3.88837097e-01,
 -4.60708593e-01, -1.39251955e-01,  2.98012847e-01,  3.79104304e-01,
  8.31154316e-02, -1.50330682e-01, -3.90226320e-02,  2.51932563e-01,
  4.71426386e-01,  5.84965643e-01,  6.08954742e-01,  4.80960066e-01,
  2.86928101e-01,  3.27027071e-01,  6.99874764e-01,  1.04476512e+00,
  9.83745392e-01,  6.54830553e-01,  5.02799063e-01,  6.61581895e-01,
  8.73326226e-01,  9.50613188e-01,  9.59502583e-01,  9.37320940e-01,
  7.96564634e-01,  6.04379740e-01,  6.18708692e-01,  8.80247202e-01,
  1.05791100e+00,  9.08379059e-01,  6.41152443e-01,  5.85284766e-01,
  7.10988232e-01,  7.70196831e-01,  7.38455424e-01,  7.77429779e-01,
  8.58005405e-01,  7.88372951e-01,  6.06711342e-01,  5.88511583e-01,
  7.99724820e-01,  9.70331048e-01,  9.24220136e-01,  8.28605155e-01,
  8.59685419e-01,  9.13774693e-01,  8.69175602e-01,  8.72188609e-01,
  1.07453927e+00,  1.28424429e+00,  1.21247454e+00,  9.53548546e-01,
  8.75435056e-01,  1.07634364e+00,  1.28534206e+00,  1.30918215e+00,
  1.24309389e+00,  1.18125090e+00,  1.05949031e+00,  9.13919870e-01,
  9.67364880e-01,  1.24814613e+00,  1.40082346e+00,  1.14809907e+00,
  7.34094247e-01,  6.09259864e-01,  8.20143780e-01,  1.02323945e+00,
  1.00446627e+00,  8.52731846e-01,  6.67398308e-01,  4.52640557e-01,
  3.28310509e-01,  4.80969629e-01,  7.90644523e-01,  8.38559722e-01,
  4.71336163e-01,  7.84638352e-02,  8.27776741e-02,  3.88569424e-01,
  5.92417691e-01,  5.43002347e-01,  3.93217627e-01,  2.49844953e-01,
  1.16819473e-01,  1.07395934e-01,  3.43268774e-01,  6.32875853e-01,
  6.06098622e-01,  2.52231762e-01,  5.75314437e-04,  1.34446852e-01,
  4.23311521e-01,  5.13071324e-01,  4.01307753e-01,  2.89347294e-01,
  2.07938839e-01,  9.07599716e-02,  4.18117043e-02,  1.87252547e-01,
  3.55531490e-01,  2.52568797e-01, -6.89479989e-02, -2.50676173e-01,
 -1.61877825e-01, -5.85027205e-02, -1.35414235e-01, -2.56642072e-01,
 -2.79535555e-01, -3.29581548e-01, -5.24048182e-01, -6.84627435e-01,
 -6.10939127e-01, -4.51121919e-01, -4.92080114e-01, -7.08300294e-01,
 -8.36091211e-01, -8.14085305e-01, -8.14025989e-01, -8.64133163e-01,
 -8.02190796e-01, -6.50167502e-01, -6.74384487e-01, -9.37081873e-01,
 -1.11121374e+00, -9.45707298e-01, -6.49586060e-01, -5.72136774e-01,
 -7.18410645e-01, -8.50289134e-01, -8.86833971e-01, -8.97476393e-01,
 -8.32938424e-01, -6.14383124e-01, -4.30629600e-01, -5.74468760e-01,
 -9.52076594e-01, -1.10945453e+00, -8.51744912e-01, -5.19685325e-01,
 -4.98526748e-01, -7.38957186e-01, -9.58844164e-01, -1.05493215e+00,
 -1.06516704e+00, -9.51458563e-01, -7.31255025e-01, -6.64635921e-01,
 -9.60279354e-01, -1.37021710e+00, -1.42942810e+00, -1.09541433e+00,
 -8.12629504e-01, -8.93643589e-01, -1.16538930e+00, -1.32853818e+00,
 -1.34156168e+00, -1.28010108e+00, -1.11907055e+00, -8.98755113e-01
 };

// `define FILTERS_BACKPREASSURE_TEST
// `define FFT_BACKPREASSURE_TEST
real coefs_b[] = {0.00257643, 0.01030574, 0.01545861, 0.01030574, 0.00257643};
real coefs_a[] = {2.63862774,  -2.76930979, 1.33928076,  -0.24982167};
// real coefs_b[] = {1.0, 1.0, 1.0, 1.0, 1.0};
// real coefs_a[] = {-1.0,  -1.0, -1.0,  -1.0};
